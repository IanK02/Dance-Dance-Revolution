module DE1_SoC (CLOCK_50, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, KEY, LEDR, GPIO_1, SW);
    input logic CLOCK_50;// 50MHz clock.
    output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
    output logic [9:0] LEDR;
	 output logic [35:0] GPIO_1;
    input logic [3:0] KEY;// True when not pressed, False when pressed
    input logic [9:0] SW;
	 

    // Generate clk off of CLOCK_50, whichClock picks rate.
    logic [31:0] div_clk;
    parameter whichClock = 14;// not many Hz clock
	 assign reset = SW[0]; //assign reset key

    clock_divider cdiv (
        .clock(CLOCK_50),
        .reset(reset),
        .divided_clocks(div_clk)
    );

    // Clock selection; allows for easy switching between simulation and board clocks
    logic clkSelect;
    // Uncomment ONE of the following two lines depending on intention
    //assign clkSelect = CLOCK_50;           // for simulation
    assign clkSelect = div_clk[whichClock];  // for board
	 
	 //logic [9:0] lsfr_num; //number generated by the lsfr
	 logic [15:0][15:0] red_pxls; //declare the 16x16 array of red pixels
	 logic [15:0][15:0] grn_pxls; //declare the 16x16 array of green pixels
	 logic [63:0] user_presses;
	 logic [3:0] lights_lost, empty_presses;
	 
	 //set red_pxls and grn_pxls to all 0 
	 initial begin
		HEX5 = 7'b1111111;
		HEX4 = 7'b1111111;
		HEX3 = 7'b1111111;
		for(int i = 0; i < 16; i++) begin
			grn_pxls[i] = '0;
			red_pxls[i] = '0;
		end
	 end
	 //------------------------------------------------
	 //keypress logic so ensure only positive edges of the user press are counted
	 logic user_press_A, user_press_B, user_press_C, user_press_D;
	 user_in uin_A (user_press_A, clkSelect, ~KEY[0]);
	 user_in uin_B (user_press_B, clkSelect, ~KEY[1]);
	 user_in uin_C (user_press_C, clkSelect, ~KEY[2]);
	 user_in uin_D (user_press_D, clkSelect, ~KEY[3]);
	 //---------------------------------------------------------------------------
	 //logic to generate pseudo random numbers with lsfr, to be used to randomly spawn lights
	 logic [12:0] lsfrA, lsfrB, lsfrC, lsfrD;
	 //logic [12:0] randomA, randomB, randomC, randomD;
	 ten_bit_lsfr #(.START_NUM(17'b01110001111100011)) lsfr_A (lsfrA, clkSelect, reset);
	 ten_bit_lsfr #(.START_NUM(17'b11000111000001000)) lsfr_B (lsfrB, clkSelect, reset);
	 ten_bit_lsfr #(.START_NUM(17'b00111111000111111)) lsfr_C (lsfrC, clkSelect, reset);
	 ten_bit_lsfr #(.START_NUM(17'b01110111000000001)) lsfr_D (lsfrD, clkSelect, reset);
	 //---------------------------------------------------------------------------
	 //logic to randomly spawn lights as well as allow the user to adjust light spawn rate
	 logic spawnA, spawnB, spawnC, spawnD;
	 column spawn_A (spawnA, SW[9:7], clkSelect, reset, lsfrA);
	 column spawn_b (spawnB, SW[9:7], clkSelect, reset, lsfrB);
	 column spawn_C (spawnC, SW[9:7], clkSelect, reset, lsfrC);
	 column spawn_D (spawnD, SW[9:7], clkSelect, reset, lsfrD);
	 //---------------------------------------------------------------------------
	 
	 //still need to implement random light spawning as well as score tallying, everything seems to
	 //be working fine until now
		
	 light_column columnA (.pixls('{
									red_pxls[0][3:0],
									red_pxls[1][3:0],
									red_pxls[2][3:0],
									red_pxls[3][3:0],
									red_pxls[4][3:0],
									red_pxls[5][3:0],
									red_pxls[6][3:0],
									red_pxls[7][3:0],
									red_pxls[8][3:0],
									red_pxls[9][3:0],
									red_pxls[10][3:0],
									red_pxls[11][3:0],
									red_pxls[12][3:0],
									red_pxls[13][3:0],
									red_pxls[14][3:0],
									red_pxls[15][3:0]
									}), 
									.user_press(user_presses[15:0]), 
									.light_lost(lights_lost[0]), 
									.empty_press(empty_presses[0]), 
									.root_spawn_signal(spawnA),
									.user_button(user_press_A),
									.light_speed(~SW[6:3]),
									.clk(clkSelect), 
									.reset(reset));
										
	 light_column columnB (.pixls('{
									grn_pxls[0][7:4],
									grn_pxls[1][7:4],
									grn_pxls[2][7:4],
									grn_pxls[3][7:4],
									grn_pxls[4][7:4],
									grn_pxls[5][7:4],
									grn_pxls[6][7:4],
									grn_pxls[7][7:4],
									grn_pxls[8][7:4],
									grn_pxls[9][7:4],
									grn_pxls[10][7:4],
									grn_pxls[11][7:4],
									grn_pxls[12][7:4],
									grn_pxls[13][7:4],
									grn_pxls[14][7:4],
									grn_pxls[15][7:4]									
									}), 
									.user_press(user_presses[31:16]), 
									.light_lost(lights_lost[1]), 
									.empty_press(empty_presses[1]), 
									.root_spawn_signal(spawnB),
									.user_button(user_press_B),
									.light_speed(~SW[6:3]),
									.clk(clkSelect), 
									.reset(reset));
										
	 light_column columnC (.pixls({
									red_pxls[0][11:8],
									red_pxls[1][11:8],
									red_pxls[2][11:8],
									red_pxls[3][11:8],
									red_pxls[4][11:8],
									red_pxls[5][11:8],
									red_pxls[6][11:8],
									red_pxls[7][11:8],
									red_pxls[8][11:8],
									red_pxls[9][11:8],
									red_pxls[10][11:8],
									red_pxls[11][11:8],
									red_pxls[12][11:8],
									red_pxls[13][11:8],
									red_pxls[14][11:8],
									red_pxls[15][11:8]
									}), 
									.user_press(user_presses[47:32]), 
									.light_lost(lights_lost[2]), 
									.empty_press(empty_presses[2]), 
									.root_spawn_signal(spawnC),
									.user_button(user_press_C),
									.light_speed(~SW[6:3]),
									.clk(clkSelect), 
									.reset(reset));
										
	 light_column columnD (.pixls({
									grn_pxls[0][15:12],
									grn_pxls[1][15:12],
									grn_pxls[2][15:12],
									grn_pxls[3][15:12],
									grn_pxls[4][15:12],
									grn_pxls[5][15:12],
									grn_pxls[6][15:12],
									grn_pxls[7][15:12],
									grn_pxls[8][15:12],
									grn_pxls[9][15:12],
									grn_pxls[10][15:12],
									grn_pxls[11][15:12],
									grn_pxls[12][15:12],
									grn_pxls[13][15:12],
									grn_pxls[14][15:12],
									grn_pxls[15][15:12]									
									}), 
									.user_press(user_presses[63:48]), 
									.light_lost(lights_lost[3]), 
									.empty_press(empty_presses[3]), 
									.root_spawn_signal(spawnD),
									.user_button(user_press_D),
									.light_speed(~SW[6:3]),
									.clk(clkSelect), 
									.reset(reset));
										
	 //score counting module
	 score_tally scoreboard (HEX0, HEX1, HEX2, user_presses, lights_lost, empty_presses, clkSelect, reset);

	 //LED Driver module 									
	 LEDDriver Driver (.CLK(clkSelect), .RST(reset), .EnableCount(1'b1), .RedPixels(red_pxls), .GrnPixels(grn_pxls), .GPIO_1);



endmodule

module DE1_SoC_testbench();
    logic CLOCK_50;
    logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
    logic [9:0] LEDR;
    logic [3:0] KEY;
    logic [9:0] SW;
	 logic [35:0] GPIO_1;

    DE1_SoC dut (CLOCK_50, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, KEY, LEDR, GPIO_1, SW);
	 
	 //assign SW[3:0] = 4'b0001;

    // Set up a simulated clock.
    parameter CLOCK_PERIOD = 100;
    initial begin
        CLOCK_50 <= 0;
        forever #(CLOCK_PERIOD/2) CLOCK_50 <= ~CLOCK_50; // Forever toggle the clock
    end
	 
	 initial begin
			SW[0] <= 1; SW[6:3] <= 4'b0000; SW[9:7] = 3'b111; @(posedge CLOCK_50); //set speed/spawning to maximum
			repeat(3) @(posedge CLOCK_50);
			SW[0] <= 0; KEY[3:0] <= 4'b1111; @(posedge CLOCK_50); //reset the machine
			//------------------------------
			repeat(5); @(posedge CLOCK_50);  //wait a bit
			//------------------------------
			//repeat(5) begin
			KEY[3] <= 0; @(posedge CLOCK_50); //user makes multiple empty presses
			KEY[3] <= 1; @(posedge CLOCK_50);
			//end
			repeat(87) @(posedge CLOCK_50);  
			KEY[3] <= 0; @(posedge CLOCK_50); //user makes winning press
			KEY[3] <= 1; @(posedge CLOCK_50);
			repeat(10) @(posedge CLOCK_50);
			KEY[1] <= 0; @(posedge CLOCK_50); //user misses
			KEY[1] <= 1; @(posedge CLOCK_50);
			repeat(16) @(posedge CLOCK_50);
			KEY[1] <= 0; @(posedge CLOCK_50); //user makes a winning press
			KEY[1] <= 1; @(posedge CLOCK_50);
			repeat(500) @(posedge CLOCK_50);
			$stop; //end simuation
	  end
endmodule